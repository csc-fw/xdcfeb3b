`timescale 1ns / 1ps

///////////////////////////////////////////////////////////////
//                                                           //
// Sub modules for DECODER                                   //
//                                                           //
///////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////
//                                                           //
// B transpose * S                                           //
//                                                           //
///////////////////////////////////////////////////////////////

module bts(
    input CLK,
    input [11:0] S,
    output reg [11:0] BTS
);

////////////////////////////////////////////////////////////////////////////////////////////////////////
// -------------------------------------------------------------------------------------------------- //
// ================================= Error Checking and Correcting code definitiions ================ //
// -------------------------------------------------------------------------------------------------- //
////////////////////////////////////////////////////////////////////////////////////////////////////////

// Rows of Parity part of Generator Matrix for ECC code Golay(24,12)
`define  BR1   12'h7FF
`define  BR2   12'hEE2
`define  BR3   12'hDC5
`define  BR4   12'hB8B
`define  BR5   12'hF16
`define  BR6   12'hE2D
`define  BR7   12'hC5B
`define  BR8   12'h8B7
`define  BR9   12'h96E
`define  BR10  12'hADC
`define  BR11  12'hDB8
`define  BR12  12'hB71


always @(posedge CLK)
begin
   BTS[11] <= ^(`BR1&S);
   BTS[10] <= ^(`BR2&S);
   BTS[9]  <= ^(`BR3&S);
   BTS[8]  <= ^(`BR4&S);
   BTS[7]  <= ^(`BR5&S);
   BTS[6]  <= ^(`BR6&S);
   BTS[5]  <= ^(`BR7&S);
   BTS[4]  <= ^(`BR8&S);
   BTS[3]  <= ^(`BR9&S);
   BTS[2]  <= ^(`BR10&S);
   BTS[1]  <= ^(`BR11&S);
   BTS[0]  <= ^(`BR12&S);
end
endmodule
